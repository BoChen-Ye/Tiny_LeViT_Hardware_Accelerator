`timescale 1ns / 1ps

package definition;
	
	parameter conv16_width=8;
	parameter conv8_width=16;
	parameter conv4_width=32;
	parameter att_width=32;
	parameter conv_Q='d1;
	parameter conv_K='d2;
	parameter conv_V='d3;
	parameter conv_att='d4;
	parameter HW=4;
endpackage
